--������ʱ����뵽����λ
--150=>2:30
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--��ʼ����
entity separatetime is
	port
	(
	clk,ce,load	: in std_logic;
	totaltime : in integer range 0 to 1440;
	ffen,sfen,fh,sh:out std_logic_vector(3 downto 0)
	);
--��������
end separatetime;
--����������one
architecture one of separatetime is
begin
--�۸�Ľ���ת��
process(clk,totaltime)
	--����һ��10λ����q
	variable comb:integer range 0 to 1441;
	variable comba,combb,combc,combd:std_logic_vector(3 downto 0);
	begin
	--��û�������ź����룬������������
	if load='0'then
		--��ʹ������Ϊ1��������������
		if ce='1' then
			--����dinΪ������ʱ��ִ���������
			if clk'event and clk='1' then
				if comb < totaltime then 
					if(comba=9 and combb=5 and combc=9)then
						comba:="0000";
						combb:="0000";
						combc:="0000";
						combd:=combd+1;
						comb:=comb+1;
					elsif(comba=9 and combb=5)then
						comba:="0000";
						combb:="0000";
						combc:=combc+1;
						comb:=comb+1;
					elsif(comba=9 and combb=5 and combc=9 and combd=5) then
						comba:="0000";
						combb:="0000";
						combc:="0000";
						combd:="0000";
						comb:=comb;
					elsif(comba=9) then
						comba:="0000";
						combb:=combb+1;
						comb:=comb+1;
					else
						comba:=comba+1;
						comb:=comb+1;
					end if;
				else
					sfen<=combb;
					ffen<=comba;
					fh<=combc;
					sh<=combd;
					comb:=totaltime;
				end if;
			end if;
		end if;	
	--�������ź�
	else
	--��ֵ����
		comb:=0;
		comba:="0000";
		combb:="0000";
		combc:="0000";
		combd:="0000";
		sfen<="0000";
		ffen<="0000";
		sh<="0000";
	end if;
	--��������
	end process;
--����������
end one;
