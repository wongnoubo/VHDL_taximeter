--�����������
--���ø���ͷ�ļ�
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--��ʼ����dp
entity total_run is
	
	port
	(
		--����ceΪ�߼����룬������ʹ�ܣ�����1��Ч���Ӹߵ����ж�ģ�����
		ce:in std_logic;
		--����clkΪ�߼����룬����������ʱ��
		clk:in std_logic;
		--����dinΪ�߼����룬���������복�����̲������ٶ�����
		din:in std_logic;
		--����dpΪ�߼����������������ж��źţ����0�����������н������1������ֹͣ
		load:in std_logic;
		--ÿ��������'1'->1km
		dp_total:out std_logic
	);
	--��������
end entity total_run;
	--����һ��������
architecture totalrun of total_run is
		--����һ���ź�dp_test������ʱ��
		--signal dp_test  : std_logic;	
	begin
		--����һ������
		process(clk,din)
		--����һ������run
		variable run : std_logic_vector(12 downto 0):="0000000000000";
		--����һ������twofive�����ź��ж�
		variable twofive : std_logic_vector(2 downto 0):=(others=>'0');
		variable twenty : std_logic_vector(3 downto 0):=(others=>'0');
			begin	
					if load='0' then
					--��ceΪ1ʱ��ִ���������
					if ce='1' then
						--��clkΪ������ʱִ���������
						if clk'event and clk='1' then
							if din='1' then
								--����500m
								if run < 250 then
									run:=run+1;
									dp_total<='0';
								else
									--����500m
									if run=250 then
										twofive:=twofive+1;
									end if;
									if run<500 then
										run:=run+1;
										dp_total<='0';
									else
										twofive:=twofive+1;
										dp_total<='1';
										twenty:=twenty+1;
										run:="0000000000000";
									end if;
								end if;
							end if;
						end if;
					end if;
				else
					run:="0000000000000";
					twofive:=(others=>'0');
					twenty:=(others=>'0');
					dp_total<='0';
				end if;
			--��������
			end process;
	--����������
	end architecture totalrun;
