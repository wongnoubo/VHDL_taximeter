--��������
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--��������
entity remove_jitter is
	port
	(
		--����ceΪ�߼����룬��Ϊʹ�ܣ�����1��Ч
		ce	: in std_logic;
		--����clkΪ�߼����룬��Ϊ��������
		clk	: in std_logic;
		--����loadΪ�߼����룬��Ϊ�����ź�
		load : in std_logic;
		--�������룬ÿ��ֻ��һ����������
		key_in	: in std_logic;
		--������İ����ź�
		key_out	: out std_logic
	);
end remove_jitter;

architecture bhv of remove_jitter is
	--��ﵽ����ʱ������
	signal N : integer := 2;
	--������
	signal count : integer range 0 to 9;
begin
	process ( clk , key_in )
	begin
		if ( clk'event and clk = '1')
		then
			--�а�������
			if ( key_in = '1' )
			then
				--ѭ��,�������������������
				if ( count = N )
				then 
					count <= count ;
				else 
					count <= count + 1;
				end if;
				--�����������������ڣ����жϰ���
				if ( count = N - 1)
				then
					key_out <= '0';
				else 
					key_out <= '1';
				end if;
			else 
				count <= 0;
			end if;
		end if;
	end process;
end bhv;
				