--���ø���ͷ�ļ�
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--��ʼ����dp
entity licheng is
	
	port
	(
		--����ceΪ�߼����룬������ʹ�ܣ�����1��Ч���Ӹߵ����ж�ģ�����
		ce:in std_logic;
		--����clkΪ�߼����룬����������ʱ��
		clk:in std_logic;
		--����dinΪ�߼����룬���������복�����̲������ٶ�����
		din:in std_logic;
		--����dpΪ�߼����������������ж��źţ����0�����������н������1������ֹͣ
		load:in std_logic;
		--�ߵ����ж������ź�
		cein:in std_logic;
		--ÿ��������'1'->1km
		dp:out std_logic;
		--��2.5km�ж�����'0'->����2.5km;'1'->2.5km����
		qibu:out std_logic;
		--Զ��12km�ж�����'0'->����12km;'1'->12km����
		yuancheng:out std_logic
	);
	--��������
	end entity licheng;
	--����һ��������
	architecture one of licheng is
		--����һ���ź�dp_test������ʱ��
		--signal dp_test  : std_logic;	
		signal flag : integer range 0 to 1:=0;
	begin
		--����һ������
		process(clk,din,cein)
		--����һ������run
		variable run : std_logic_vector(12 downto 0):="0000000000000";
		--����һ������twofive�����ź��ж�
		variable twofive : std_logic_vector(2 downto 0):=(others=>'0');
		variable twenty : std_logic_vector(3 downto 0):=(others=>'0');
			begin	
			if load='0' then
				--��ceΪ1ʱ��ִ���������
				if ce='1' then
					--��clkΪ������ʱִ���������
					if clk'event and clk='1' then
						if flag=0 then--��״̬����̼������ܵ��ߵ���״̬��Ӱ��
							if din='1' then
								--����500m
								if run < 250 then
									run:=run+1;
									dp<='0';
								else
									--����500m
									if run=250 then
										twofive:=twofive+1;
									end if;
									if run<500 then--
										run:=run+1;
										dp<='0';
									else
										twofive:=twofive+1;
										dp<='1';
										twenty:=twenty+1;
										run:="0000000000000";
									end if;
								end if;
							end if;
							if twenty < 12 then
								yuancheng<='0';
							else
								yuancheng<='1';
								--13
								twenty:="1101";
							end if;
							--�ж��Ƿ񵽴������
							if twofive < 4 then
								qibu<='0';
							else
								qibu<='1';
								flag<=1;
								dp<='1';
								--5
								twofive:="101";
							end if;
						end if;
						if cein='1' and flag=1 then--����״̬�½�����̼Ƽ�
							if din='1' then
								--����500m
								if run < 250 then
									run:=run+1;
									dp<='0';
								else
									--����500m
									if run=250 then
										twofive:=twofive+1;
									end if;
									if run<500 then
										run:=run+1;
										dp<='0';
									else
										twofive:=twofive+1;
										dp<='1';
										twenty:=twenty+1;
										run:="0000000000000";
									end if;
								end if;
							end if;
							if twenty < 12 then
								yuancheng<='0';
							else
								yuancheng<='1';
								--13
								twenty:="1101";
							end if;
							--�ж��Ƿ񵽴������
							if twofive < 4 then
								qibu<='0';
							else
								qibu<='1';
								flag<=1;
								--5
								twofive:="101";
							end if;
						end if;
					end if;
				end if;
			else
				qibu<='0';
				yuancheng<='0';
				run:="0000000000000";
				twofive:=(others=>'0');
				twenty:=(others=>'0');
				dp<='0';
				flag<=1;
			end if;
		--��������
		end process;
	--����������
	end architecture one;
