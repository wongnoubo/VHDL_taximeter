--���ø���ͷ�ļ�
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--��ʼ����
entity lingcheng is
	port
	(
	--����clkΪ�߼����룬��Ϊ��������
	clk	: in std_logic;
	--����loadΪ�߼����룬��Ϊ�����ź�
	timesel : in std_logic;--ʱ������ģʽ
	settime : in std_logic_vector(10 downto 0);
	--����ceoutΪ�߼��������Ϊ�жϽ�����
	ceout : out std_logic
	);
--��������
end lingcheng;

--����һ��������
architecture one of lingcheng is
begin
--����һ������
process(clk,settime)
	--����һ������dintest
	variable time:integer range 0 to 61;
	variable mins:std_logic_vector(10 downto 0):=(others=>'0');
	begin
	--û�������źţ�������������
	--clk���������أ�ִ���������
	if clk'event and clk='1' then 
		if timesel='1' then
			mins:=settime;
		end if;
		if time< 60 then 
			--������һ
			time:=time + 1;
		else
			time:=0;
			mins:=mins+1;
		end if;
		--6h
		if mins < 360 then
			ceout<='1';
		--23h
		elsif mins > 1380 and mins < 1441 then
			ceout<='1';
			--���Ϊ0���ú���ļ������Ȳ�Ҫ����
		elsif mins > 1440 then
			time:=0;
			mins:=(others=>'0');
			--���1���𲽼۽���������ļ�����������ʼ
		else
		--6h-23h
			ceout<='0';
		end if;
	end if;
	--��������
	end process;
--����������
end one;