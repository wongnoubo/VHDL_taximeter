--ͳ���������������ʵ�����з����ܵ�����
--���ø���ͷ�ļ�
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--��ʼ����
entity countplus is
	port
	(
	--����ceΪ�߼����룬��Ϊʹ�ܣ�����1��Ч
	ce	: in std_logic;
	--����loadΪ�߼����룬��Ϊ�����ź�
	load: in std_logic;
	--����
	din:in std_logic;
	--����ceoutΪ�߼��������Ϊ�жϽ�����
	total : out integer range 0 to 1440
	);
--��������
end countplus;

--����һ��������
architecture one of countplus is
begin
	process(ce,din) 
	variable comb:integer range 0 to 1440;
	begin
		if load='0' then
			if ce='1' then
				if din='1' and din'event then
					comb:=comb+1;
					total<=comb;
				end if;
			end if;
		else
			comb:=0;
			total<=0;
		end if;
	end process;
end one;
