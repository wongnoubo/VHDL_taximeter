	--���ø���ͷ�ļ�
	library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.std_logic_arith.all;
	--��ʼ����
	entity or2time is
		port
		(
		--����dinΪ�߼����룬����������ʱ���ź�
		--����loadΪ�߼����룬����������
		ce : in std_logic;
		timesel : in std_logic;--ʱ�����ñ�־
		ffen,sfen,fh,sh:in std_logic_vector(3 downto 0);--���⳵��ʻʱ����ʾ
		vffen,vsfen,vfh,vsh:in integer range 0 to 9; --����ʱ������
		rffen,rsfen,rfh,rsh:out std_logic_vector(3 downto 0)
		);
	--��������
	end or2time;
	--����������one
	architecture one of or2time is
	signal vffentemp,vsfentemp,vfhtemp,vshtemp:integer range 0 to 9;
	signal rffentemp,rsfentemp,rfhtemp,rshtemp:std_logic_vector(3 downto 0);
		begin 
	process(ce,ffen,sfen,fh,sh,vffen,vsfen,vfh,vsh)
		begin
		if ce='1' then
			vffentemp<=vffen;
			vsfentemp<=vsfen;
			vfhtemp<=vfh;
			vshtemp<=vsh;
			if timesel='1' then --����״̬
				rffentemp<=conv_std_logic_vector(vffentemp,4);
				rsfentemp<=conv_std_logic_vector(vsfentemp,4);
				rfhtemp<=conv_std_logic_vector(vfhtemp,4);
				rshtemp<=conv_std_logic_vector(vshtemp,4);
				rffen<=rffentemp;
				rsfen<=rsfentemp;
				rfh<=rfhtemp;
				rsh<=rshtemp;
			else
				rffen<=ffen;
				rsfen<=sfen;
				rfh<=fh;
				rsh<=sh;
			end if;
		end if;
		end process;
	--����������
	end one;
