--���ø���ͷ�ļ�
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--�𲽼��ڼƼ�
entity starting_price is
	--generic(
		--		day_starting_price : integer range 0 to 200 := 100;		--�����𲽼�
		--		night_starting_price : integer range 0 to 200 := 120		--ҹ���𲽼�
	--);
		port(
				st : in std_logic;
				load : in std_logic;
				--night drive
				night : in std_logic;
				--ʱ������
				clk : in std_logic;
				--����״̬���жϵļƼ�״̬
				state_pricing : in integer range 1 to 4;
				--����
				day_starting_price :in integer range 0 to 200;
				night_starting_price :in integer range 0 to 200;
				total_price : out integer range 0 to 10000
	);
end entity starting_price;

architecture start of starting_price is
begin
	process(load , clk ,  night , state_pricing  )
	begin
		if state_pricing = 1 and load = '1' then    --�ܼ۸�λΪ0
			total_price <= 0;
		end if;
		if state_pricing = 2 then                    --�𲽼��ڼƼ�
			if night = '0' then							--�����𲽼�
				total_price <= day_starting_price;
			elsif night = '1' then						--ҹ���𲽼�
				total_price <= night_starting_price;
			end if;
		end if;
		if state_pricing = 3 then
			total_price <= 0;
		end if;
	end process;
end start;