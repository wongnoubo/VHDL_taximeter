	--���ø���ͷ�ļ�
	library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	--��ʼ����
	entity or2total is
		port
		(
		--����dinΪ�߼����룬����������ʱ���ź�
		--����loadΪ�߼����룬����������
		ce : in std_logic;
		pricesel : in integer;--�۸�λ��ѡ��
		total1	: in integer range 0 to 9999;--�𲽼���Ƽ�
		total2	: in integer range 0 to 9999;--�𲽼��ڼƼ�
		price : in integer range 0 to 9999;--���ü۸�Ƽ�
		total	: out integer range 0 to 9999
		);
	--��������
	end or2total;
	--����������one
	architecture one of or2total is
		begin
	process(ce,total1,total2)
		begin
		if ce='1' then
			if total1>0 and total2=0 and pricesel=0 then
				total<=total1;
			elsif total1=0 and total2>0 and pricesel=0 then
				total<=total2;
			elsif pricesel>0 then
				total<=price;
			end if;
		end if;
		end process;
	--����������
	end one;
