--����Ʊ�۸��ո�ʮ��ǧ���ηֿ�
--���ø���ͷ�ļ�
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
--��ʼ����
entity separateprice is
	port
	(
	clk,ce,load	: in std_logic;
	total : in integer range 0 to 10000;
	dout : out std_logic;
	ge,shi,bai,qian,wan:out std_logic_vector(3 downto 0)
	);
--��������
end separateprice;
--����������one
architecture one of separateprice is
begin
--�۸�Ľ���ת��
process(clk,total)
	--����һ��10λ����q
	variable comb:integer range 0 to 10001;
	variable comba,combb,combc,combd,combe:std_logic_vector(3 downto 0);
	begin
	--��û�������ź����룬������������
	if load='0'then
		--��ʹ������Ϊ1��������������
		if ce='1' then
			--����dinΪ������ʱ��ִ���������
			if clk'event and clk='1' then
				if comb < total then 
					if(comba=9 and combb=9 and combc=9)then
						comba:="0000";
						combb:="0000";
						combc:="0000";
						combd:=combd+1;
						comb:=comb+1;
					elsif(comba=9 and combb=9)then
						comba:="0000";
						combb:="0000";
						combc:=combc+1;
						comb:=comb+1;
					elsif(comba=9 and combb=9 and combc=9 and combd=9) then
						comba:="0000";
						combb:="0000";
						combc:="0000";
						combd:="0000";
						combe:=combe+1;
						comb:=comb+1;
					elsif(comba=9) then
						comba:="0000";
						combb:=combb+1;
						comb:=comb+1;
					else
						comba:=comba+1;
						comb:=comb+1;
					end if;
				else
					shi<=combb;
					ge<=comba;
					bai<=combc;
					qian<=combd;
					wan<=combe;
					comb:=total;
				end if;
			end if;
		end if;	
	--�������ź�
	else
	--��ֵ����
		comb:=0;
		comba:="0000";
		combb:="0000";
		combc:="0000";
		combd:="0000";
		combe:="0000";
		shi<="0000";
		ge<="0000";
		bai<="0000";
		qian<="0000";
		wan<="0000";
	end if;
	--��������
	end process;
--����������
end one;
